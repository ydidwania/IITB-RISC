// instantiating_memory_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module instantiating_memory_system (
		input  wire        system_0_onchip_memory_0_clk1_clk,         //   system_0_onchip_memory_0_clk1.clk
		input  wire        system_0_onchip_memory_0_reset1_reset,     // system_0_onchip_memory_0_reset1.reset
		input  wire        system_0_onchip_memory_0_reset1_reset_req, //                                .reset_req
		input  wire [15:0] system_0_onchip_memory_0_s1_address,       //     system_0_onchip_memory_0_s1.address
		input  wire        system_0_onchip_memory_0_s1_clken,         //                                .clken
		input  wire        system_0_onchip_memory_0_s1_chipselect,    //                                .chipselect
		input  wire        system_0_onchip_memory_0_s1_write,         //                                .write
		output wire [15:0] system_0_onchip_memory_0_s1_readdata,      //                                .readdata
		input  wire [15:0] system_0_onchip_memory_0_s1_writedata,     //                                .writedata
		input  wire [1:0]  system_0_onchip_memory_0_s1_byteenable     //                                .byteenable
	);

	instantiating_memory_system_system_0 system_0 (
		.onchip_memory_0_clk1_clk         (system_0_onchip_memory_0_clk1_clk),         //   onchip_memory_0_clk1.clk
		.onchip_memory_0_reset1_reset     (system_0_onchip_memory_0_reset1_reset),     // onchip_memory_0_reset1.reset
		.onchip_memory_0_reset1_reset_req (system_0_onchip_memory_0_reset1_reset_req), //                       .reset_req
		.onchip_memory_0_s1_address       (system_0_onchip_memory_0_s1_address),       //     onchip_memory_0_s1.address
		.onchip_memory_0_s1_clken         (system_0_onchip_memory_0_s1_clken),         //                       .clken
		.onchip_memory_0_s1_chipselect    (system_0_onchip_memory_0_s1_chipselect),    //                       .chipselect
		.onchip_memory_0_s1_write         (system_0_onchip_memory_0_s1_write),         //                       .write
		.onchip_memory_0_s1_readdata      (system_0_onchip_memory_0_s1_readdata),      //                       .readdata
		.onchip_memory_0_s1_writedata     (system_0_onchip_memory_0_s1_writedata),     //                       .writedata
		.onchip_memory_0_s1_byteenable    (system_0_onchip_memory_0_s1_byteenable)     //                       .byteenable
	);

endmodule
