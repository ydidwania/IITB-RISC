// instantiating_memory_system_system_0.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module instantiating_memory_system_system_0 (
		input  wire        onchip_memory_0_clk1_clk,         //   onchip_memory_0_clk1.clk
		input  wire        onchip_memory_0_reset1_reset,     // onchip_memory_0_reset1.reset
		input  wire        onchip_memory_0_reset1_reset_req, //                       .reset_req
		input  wire [15:0] onchip_memory_0_s1_address,       //     onchip_memory_0_s1.address
		input  wire        onchip_memory_0_s1_clken,         //                       .clken
		input  wire        onchip_memory_0_s1_chipselect,    //                       .chipselect
		input  wire        onchip_memory_0_s1_write,         //                       .write
		output wire [15:0] onchip_memory_0_s1_readdata,      //                       .readdata
		input  wire [15:0] onchip_memory_0_s1_writedata,     //                       .writedata
		input  wire [1:0]  onchip_memory_0_s1_byteenable     //                       .byteenable
	);

	instantiating_memory_system_system_0_onchip_memory_0 onchip_memory_0 (
		.clk        (onchip_memory_0_clk1_clk),         //   clk1.clk
		.address    (onchip_memory_0_s1_address),       //     s1.address
		.clken      (onchip_memory_0_s1_clken),         //       .clken
		.chipselect (onchip_memory_0_s1_chipselect),    //       .chipselect
		.write      (onchip_memory_0_s1_write),         //       .write
		.readdata   (onchip_memory_0_s1_readdata),      //       .readdata
		.writedata  (onchip_memory_0_s1_writedata),     //       .writedata
		.byteenable (onchip_memory_0_s1_byteenable),    //       .byteenable
		.reset      (onchip_memory_0_reset1_reset),     // reset1.reset
		.reset_req  (onchip_memory_0_reset1_reset_req), //       .reset_req
		.freeze     (1'b0)                              // (terminated)
	);

endmodule
