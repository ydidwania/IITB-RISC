library ieee;	
use ieee.std_logic_1164.all;

entity mux3bit2to1 is
	port(in_1,in_2       : in std_logic_vector(0 to 2);
		sel 	     : in std_logic;
		mux_out	     : out std_logic_vector(0 to 2));
end entity;

architecture behave of mux3bit2to1 is
begin
	process(sel)
	begin
		case sel is
		when '0' =>
			mux_out <= in_1;
		when '1' =>
			mux_out <= in_2;
		end case;
	end process;
end behave;
